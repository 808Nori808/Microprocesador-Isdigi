hola soy hugo